--------------------------------------------------------------------------------
--                       FixFunctionByTable_Freq1_uid2
-- Evaluator for log(x+0.1)/log(2) on [0,1) for lsbIn=-9 (wIn=9), msbout=2, lsbOut=-3 (wOut=6). Out interval: [-3.32193; 0.13494]. Output is signed

-- VHDL generated for Kintex7 @ 1MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2010-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1000
-- Target frequency (MHz): 1
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: Y: (c0, 0.543000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixFunctionByTable_Freq1_uid2 is
    port (X : in  std_logic_vector(8 downto 0);
          Y : out  std_logic_vector(5 downto 0)   );
end entity;

architecture arch of FixFunctionByTable_Freq1_uid2 is
signal Y0 :  std_logic_vector(5 downto 0);
   -- timing of Y0: (c0, 0.543000ns)
signal Y1 :  std_logic_vector(5 downto 0);
   -- timing of Y1: (c0, 0.543000ns)
begin
   with X  select  Y0 <= 
      "100101" when "000000000",
      "100110" when "000000001",
      "100110" when "000000010",
      "100110" when "000000011",
      "100110" when "000000100",
      "100110" when "000000101",
      "100111" when "000000110",
      "100111" when "000000111",
      "100111" when "000001000",
      "100111" when "000001001",
      "100111" when "000001010",
      "101000" when "000001011",
      "101000" when "000001100",
      "101000" when "000001101",
      "101000" when "000001110",
      "101000" when "000001111",
      "101001" when "000010000",
      "101001" when "000010001",
      "101001" when "000010010",
      "101001" when "000010011",
      "101001" when "000010100",
      "101001" when "000010101",
      "101010" when "000010110",
      "101010" when "000010111",
      "101010" when "000011000",
      "101010" when "000011001",
      "101010" when "000011010",
      "101010" when "000011011",
      "101010" when "000011100",
      "101011" when "000011101",
      "101011" when "000011110",
      "101011" when "000011111",
      "101011" when "000100000",
      "101011" when "000100001",
      "101011" when "000100010",
      "101011" when "000100011",
      "101100" when "000100100",
      "101100" when "000100101",
      "101100" when "000100110",
      "101100" when "000100111",
      "101100" when "000101000",
      "101100" when "000101001",
      "101100" when "000101010",
      "101100" when "000101011",
      "101101" when "000101100",
      "101101" when "000101101",
      "101101" when "000101110",
      "101101" when "000101111",
      "101101" when "000110000",
      "101101" when "000110001",
      "101101" when "000110010",
      "101101" when "000110011",
      "101110" when "000110100",
      "101110" when "000110101",
      "101110" when "000110110",
      "101110" when "000110111",
      "101110" when "000111000",
      "101110" when "000111001",
      "101110" when "000111010",
      "101110" when "000111011",
      "101110" when "000111100",
      "101110" when "000111101",
      "101111" when "000111110",
      "101111" when "000111111",
      "101111" when "001000000",
      "101111" when "001000001",
      "101111" when "001000010",
      "101111" when "001000011",
      "101111" when "001000100",
      "101111" when "001000101",
      "101111" when "001000110",
      "101111" when "001000111",
      "110000" when "001001000",
      "110000" when "001001001",
      "110000" when "001001010",
      "110000" when "001001011",
      "110000" when "001001100",
      "110000" when "001001101",
      "110000" when "001001110",
      "110000" when "001001111",
      "110000" when "001010000",
      "110000" when "001010001",
      "110000" when "001010010",
      "110001" when "001010011",
      "110001" when "001010100",
      "110001" when "001010101",
      "110001" when "001010110",
      "110001" when "001010111",
      "110001" when "001011000",
      "110001" when "001011001",
      "110001" when "001011010",
      "110001" when "001011011",
      "110001" when "001011100",
      "110001" when "001011101",
      "110001" when "001011110",
      "110010" when "001011111",
      "110010" when "001100000",
      "110010" when "001100001",
      "110010" when "001100010",
      "110010" when "001100011",
      "110010" when "001100100",
      "110010" when "001100101",
      "110010" when "001100110",
      "110010" when "001100111",
      "110010" when "001101000",
      "110010" when "001101001",
      "110010" when "001101010",
      "110010" when "001101011",
      "110011" when "001101100",
      "110011" when "001101101",
      "110011" when "001101110",
      "110011" when "001101111",
      "110011" when "001110000",
      "110011" when "001110001",
      "110011" when "001110010",
      "110011" when "001110011",
      "110011" when "001110100",
      "110011" when "001110101",
      "110011" when "001110110",
      "110011" when "001110111",
      "110011" when "001111000",
      "110011" when "001111001",
      "110011" when "001111010",
      "110100" when "001111011",
      "110100" when "001111100",
      "110100" when "001111101",
      "110100" when "001111110",
      "110100" when "001111111",
      "110100" when "010000000",
      "110100" when "010000001",
      "110100" when "010000010",
      "110100" when "010000011",
      "110100" when "010000100",
      "110100" when "010000101",
      "110100" when "010000110",
      "110100" when "010000111",
      "110100" when "010001000",
      "110100" when "010001001",
      "110101" when "010001010",
      "110101" when "010001011",
      "110101" when "010001100",
      "110101" when "010001101",
      "110101" when "010001110",
      "110101" when "010001111",
      "110101" when "010010000",
      "110101" when "010010001",
      "110101" when "010010010",
      "110101" when "010010011",
      "110101" when "010010100",
      "110101" when "010010101",
      "110101" when "010010110",
      "110101" when "010010111",
      "110101" when "010011000",
      "110101" when "010011001",
      "110101" when "010011010",
      "110110" when "010011011",
      "110110" when "010011100",
      "110110" when "010011101",
      "110110" when "010011110",
      "110110" when "010011111",
      "110110" when "010100000",
      "110110" when "010100001",
      "110110" when "010100010",
      "110110" when "010100011",
      "110110" when "010100100",
      "110110" when "010100101",
      "110110" when "010100110",
      "110110" when "010100111",
      "110110" when "010101000",
      "110110" when "010101001",
      "110110" when "010101010",
      "110110" when "010101011",
      "110110" when "010101100",
      "110110" when "010101101",
      "110111" when "010101110",
      "110111" when "010101111",
      "110111" when "010110000",
      "110111" when "010110001",
      "110111" when "010110010",
      "110111" when "010110011",
      "110111" when "010110100",
      "110111" when "010110101",
      "110111" when "010110110",
      "110111" when "010110111",
      "110111" when "010111000",
      "110111" when "010111001",
      "110111" when "010111010",
      "110111" when "010111011",
      "110111" when "010111100",
      "110111" when "010111101",
      "110111" when "010111110",
      "110111" when "010111111",
      "110111" when "011000000",
      "110111" when "011000001",
      "111000" when "011000010",
      "111000" when "011000011",
      "111000" when "011000100",
      "111000" when "011000101",
      "111000" when "011000110",
      "111000" when "011000111",
      "111000" when "011001000",
      "111000" when "011001001",
      "111000" when "011001010",
      "111000" when "011001011",
      "111000" when "011001100",
      "111000" when "011001101",
      "111000" when "011001110",
      "111000" when "011001111",
      "111000" when "011010000",
      "111000" when "011010001",
      "111000" when "011010010",
      "111000" when "011010011",
      "111000" when "011010100",
      "111000" when "011010101",
      "111000" when "011010110",
      "111000" when "011010111",
      "111000" when "011011000",
      "111001" when "011011001",
      "111001" when "011011010",
      "111001" when "011011011",
      "111001" when "011011100",
      "111001" when "011011101",
      "111001" when "011011110",
      "111001" when "011011111",
      "111001" when "011100000",
      "111001" when "011100001",
      "111001" when "011100010",
      "111001" when "011100011",
      "111001" when "011100100",
      "111001" when "011100101",
      "111001" when "011100110",
      "111001" when "011100111",
      "111001" when "011101000",
      "111001" when "011101001",
      "111001" when "011101010",
      "111001" when "011101011",
      "111001" when "011101100",
      "111001" when "011101101",
      "111001" when "011101110",
      "111001" when "011101111",
      "111001" when "011110000",
      "111010" when "011110001",
      "111010" when "011110010",
      "111010" when "011110011",
      "111010" when "011110100",
      "111010" when "011110101",
      "111010" when "011110110",
      "111010" when "011110111",
      "111010" when "011111000",
      "111010" when "011111001",
      "111010" when "011111010",
      "111010" when "011111011",
      "111010" when "011111100",
      "111010" when "011111101",
      "111010" when "011111110",
      "111010" when "011111111",
      "111010" when "100000000",
      "111010" when "100000001",
      "111010" when "100000010",
      "111010" when "100000011",
      "111010" when "100000100",
      "111010" when "100000101",
      "111010" when "100000110",
      "111010" when "100000111",
      "111010" when "100001000",
      "111010" when "100001001",
      "111010" when "100001010",
      "111011" when "100001011",
      "111011" when "100001100",
      "111011" when "100001101",
      "111011" when "100001110",
      "111011" when "100001111",
      "111011" when "100010000",
      "111011" when "100010001",
      "111011" when "100010010",
      "111011" when "100010011",
      "111011" when "100010100",
      "111011" when "100010101",
      "111011" when "100010110",
      "111011" when "100010111",
      "111011" when "100011000",
      "111011" when "100011001",
      "111011" when "100011010",
      "111011" when "100011011",
      "111011" when "100011100",
      "111011" when "100011101",
      "111011" when "100011110",
      "111011" when "100011111",
      "111011" when "100100000",
      "111011" when "100100001",
      "111011" when "100100010",
      "111011" when "100100011",
      "111011" when "100100100",
      "111011" when "100100101",
      "111011" when "100100110",
      "111011" when "100100111",
      "111100" when "100101000",
      "111100" when "100101001",
      "111100" when "100101010",
      "111100" when "100101011",
      "111100" when "100101100",
      "111100" when "100101101",
      "111100" when "100101110",
      "111100" when "100101111",
      "111100" when "100110000",
      "111100" when "100110001",
      "111100" when "100110010",
      "111100" when "100110011",
      "111100" when "100110100",
      "111100" when "100110101",
      "111100" when "100110110",
      "111100" when "100110111",
      "111100" when "100111000",
      "111100" when "100111001",
      "111100" when "100111010",
      "111100" when "100111011",
      "111100" when "100111100",
      "111100" when "100111101",
      "111100" when "100111110",
      "111100" when "100111111",
      "111100" when "101000000",
      "111100" when "101000001",
      "111100" when "101000010",
      "111100" when "101000011",
      "111100" when "101000100",
      "111100" when "101000101",
      "111100" when "101000110",
      "111101" when "101000111",
      "111101" when "101001000",
      "111101" when "101001001",
      "111101" when "101001010",
      "111101" when "101001011",
      "111101" when "101001100",
      "111101" when "101001101",
      "111101" when "101001110",
      "111101" when "101001111",
      "111101" when "101010000",
      "111101" when "101010001",
      "111101" when "101010010",
      "111101" when "101010011",
      "111101" when "101010100",
      "111101" when "101010101",
      "111101" when "101010110",
      "111101" when "101010111",
      "111101" when "101011000",
      "111101" when "101011001",
      "111101" when "101011010",
      "111101" when "101011011",
      "111101" when "101011100",
      "111101" when "101011101",
      "111101" when "101011110",
      "111101" when "101011111",
      "111101" when "101100000",
      "111101" when "101100001",
      "111101" when "101100010",
      "111101" when "101100011",
      "111101" when "101100100",
      "111101" when "101100101",
      "111101" when "101100110",
      "111101" when "101100111",
      "111101" when "101101000",
      "111101" when "101101001",
      "111110" when "101101010",
      "111110" when "101101011",
      "111110" when "101101100",
      "111110" when "101101101",
      "111110" when "101101110",
      "111110" when "101101111",
      "111110" when "101110000",
      "111110" when "101110001",
      "111110" when "101110010",
      "111110" when "101110011",
      "111110" when "101110100",
      "111110" when "101110101",
      "111110" when "101110110",
      "111110" when "101110111",
      "111110" when "101111000",
      "111110" when "101111001",
      "111110" when "101111010",
      "111110" when "101111011",
      "111110" when "101111100",
      "111110" when "101111101",
      "111110" when "101111110",
      "111110" when "101111111",
      "111110" when "110000000",
      "111110" when "110000001",
      "111110" when "110000010",
      "111110" when "110000011",
      "111110" when "110000100",
      "111110" when "110000101",
      "111110" when "110000110",
      "111110" when "110000111",
      "111110" when "110001000",
      "111110" when "110001001",
      "111110" when "110001010",
      "111110" when "110001011",
      "111110" when "110001100",
      "111110" when "110001101",
      "111110" when "110001110",
      "111111" when "110001111",
      "111111" when "110010000",
      "111111" when "110010001",
      "111111" when "110010010",
      "111111" when "110010011",
      "111111" when "110010100",
      "111111" when "110010101",
      "111111" when "110010110",
      "111111" when "110010111",
      "111111" when "110011000",
      "111111" when "110011001",
      "111111" when "110011010",
      "111111" when "110011011",
      "111111" when "110011100",
      "111111" when "110011101",
      "111111" when "110011110",
      "111111" when "110011111",
      "111111" when "110100000",
      "111111" when "110100001",
      "111111" when "110100010",
      "111111" when "110100011",
      "111111" when "110100100",
      "111111" when "110100101",
      "111111" when "110100110",
      "111111" when "110100111",
      "111111" when "110101000",
      "111111" when "110101001",
      "111111" when "110101010",
      "111111" when "110101011",
      "111111" when "110101100",
      "111111" when "110101101",
      "111111" when "110101110",
      "111111" when "110101111",
      "111111" when "110110000",
      "111111" when "110110001",
      "111111" when "110110010",
      "111111" when "110110011",
      "111111" when "110110100",
      "111111" when "110110101",
      "111111" when "110110110",
      "111111" when "110110111",
      "000000" when "110111000",
      "000000" when "110111001",
      "000000" when "110111010",
      "000000" when "110111011",
      "000000" when "110111100",
      "000000" when "110111101",
      "000000" when "110111110",
      "000000" when "110111111",
      "000000" when "111000000",
      "000000" when "111000001",
      "000000" when "111000010",
      "000000" when "111000011",
      "000000" when "111000100",
      "000000" when "111000101",
      "000000" when "111000110",
      "000000" when "111000111",
      "000000" when "111001000",
      "000000" when "111001001",
      "000000" when "111001010",
      "000000" when "111001011",
      "000000" when "111001100",
      "000000" when "111001101",
      "000000" when "111001110",
      "000000" when "111001111",
      "000000" when "111010000",
      "000000" when "111010001",
      "000000" when "111010010",
      "000000" when "111010011",
      "000000" when "111010100",
      "000000" when "111010101",
      "000000" when "111010110",
      "000000" when "111010111",
      "000000" when "111011000",
      "000000" when "111011001",
      "000000" when "111011010",
      "000000" when "111011011",
      "000000" when "111011100",
      "000000" when "111011101",
      "000000" when "111011110",
      "000000" when "111011111",
      "000000" when "111100000",
      "000000" when "111100001",
      "000000" when "111100010",
      "000000" when "111100011",
      "000001" when "111100100",
      "000001" when "111100101",
      "000001" when "111100110",
      "000001" when "111100111",
      "000001" when "111101000",
      "000001" when "111101001",
      "000001" when "111101010",
      "000001" when "111101011",
      "000001" when "111101100",
      "000001" when "111101101",
      "000001" when "111101110",
      "000001" when "111101111",
      "000001" when "111110000",
      "000001" when "111110001",
      "000001" when "111110010",
      "000001" when "111110011",
      "000001" when "111110100",
      "000001" when "111110101",
      "000001" when "111110110",
      "000001" when "111110111",
      "000001" when "111111000",
      "000001" when "111111001",
      "000001" when "111111010",
      "000001" when "111111011",
      "000001" when "111111100",
      "000001" when "111111101",
      "000001" when "111111110",
      "000001" when "111111111",
      "------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

